../../../TheSDK_generators/verilog/f2_tx_dsp.v