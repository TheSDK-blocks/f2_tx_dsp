../../../TheSDK_generators/verilog/tb_f2_tx_dsp.v